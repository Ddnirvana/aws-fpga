module test (
clk,
test_input,
test_output,
test_inout
);

inout clk;
input test_input;
output test_output;
inout test_inout;

endmodule