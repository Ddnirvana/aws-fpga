module test (
clk,
test_input
);

input clk;
input test_input;

endmodule