module test (
clk,
test1
);

input clk;
inout test1;

endmodule