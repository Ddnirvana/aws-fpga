module test (
clk,
test_input,
test_output,
test_inout
);

input clk;
input test_input;
output test_output;
inout test_inout;

wire clk;
wire test_input;
wire test_output;
wire test_inout;

endmodule