module test (
clk,
test1
);

input clk;
input test1;

endmodule