module test (
clk,
test_input,
test_output
);

input clk;
input test_input;
output test_output;

endmodule